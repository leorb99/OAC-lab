/*`ifndef PARAM
	`include "Parametros.v"
`endif

module Control ()*/